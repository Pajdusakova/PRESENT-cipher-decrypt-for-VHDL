library IEEE;
use IEEE.std_logic_1164.all;

entity pLayer_dec is
	port( X: in std_logic_vector(63 downto 0);
			Y: out std_logic_vector(63 downto 0));
end pLayer_dec;

architecture rtl of pLayer_dec is
begin
	Y(63)<=X(63); Y(62)<=X(47); Y(61)<=X(31); Y(60)<=X(15);
	Y(59)<=X(62); Y(58)<=X(46); Y(57)<=X(30); Y(56)<=X(14);
	Y(55)<=X(61); Y(54)<=X(45); Y(53)<=X(29); Y(52)<=X(13);
	Y(51)<=X(60); Y(50)<=X(44); Y(49)<=X(28); Y(48)<=X(12);
	Y(47)<=X(59); Y(46)<=X(43); Y(45)<=X(27); Y(44)<=X(11);
	Y(43)<=X(58); Y(42)<=X(42); Y(41)<=X(26); Y(40)<=X(10);
	Y(39)<=X(57); Y(38)<=X(41); Y(37)<=X(25); Y(36)<=X( 9);
	Y(35)<=X(56); Y(34)<=X(40); Y(33)<=X(24); Y(32)<=X( 8);
	Y(31)<=X(55); Y(30)<=X(39); Y(29)<=X(23); Y(28)<=X( 7);
	Y(27)<=X(54); Y(26)<=X(38); Y(25)<=X(22); Y(24)<=X( 6);
	Y(23)<=X(53); Y(22)<=X(37); Y(21)<=X(21); Y(20)<=X( 5);
	Y(19)<=X(52); Y(18)<=X(36); Y(17)<=X(20); Y(16)<=X( 4);
	Y(15)<=X(51); Y(14)<=X(35); Y(13)<=X(19); Y(12)<=X( 3);
	Y(11)<=X(50); Y(10)<=X(34); Y( 9)<=X(18); Y( 8)<=X( 2);
	Y( 7)<=X(49); Y( 6)<=X(33); Y( 5)<=X(17); Y( 4)<=X( 1);
	Y( 3)<=X(48); Y( 2)<=X(32); Y( 1)<=X(16); Y( 0)<=X( 0);
end rtl;